module Average(clk, reset, data, valid, out);
input        clk, reset;
input  [7:0] data;
output       valid;
output [7:0] out;
//===================== Your Design =====================

//===================== Your Design =====================
endmodule
